module logger 

